module accumulator #(parameter INPUT_NUM=16; parameter WIDTH = 5;) ();
    output  [WIDTH-1:0] out;
    input   clk;
    input   [INPUT_NUM-1:0] in;

    // implement a tree adder



endmodule