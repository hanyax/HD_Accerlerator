

module accelerator_top #(parameter WIDTH=16) () 
    input logic clk;
    input logic [WIDTH-1:0] projection_matrix; // P matrix is binary
    
    

endmodule 